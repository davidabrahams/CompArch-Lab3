module cpuRunner;


endmodule
